module T05_port_2 (
    input wire clk,
    input pertama,
    input kedua,
    inout [15:0] data,
    output keluaran);
    
endmodule
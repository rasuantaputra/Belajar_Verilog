module T20_2_repeat;

    initial begin
        repeat (5) begin
            $display("ini iterasi menggunakan repeat loop...");
        end 
    end
    
endmodule
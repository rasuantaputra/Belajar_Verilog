// design top level

module mod3 ();
    
endmodule

module mod4 ();
    
endmodule

module mod1 ();
    
endmodule

module mod2 ();
    
endmodule

// top-level module
module T04_module3 ();
    
    wire net;

    mod1
    mod2
    
endmodule
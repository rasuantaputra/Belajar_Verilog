module T36_math_function 
#(parameter NUM_UNITS = 7)
(input [$clog2(NUM_UNITS - 1:0)] activate_unit);
    
endmodule